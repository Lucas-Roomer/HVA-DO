library ieee;
use ieee.std_logic_1164.all;

entity opdracht_231 is
	port(
		d : in std_logic;
		clk : in std_logic;
		q : out std_logic);
end entity opdracht_231;

architecture behaviour of opdracht_231 is
begin


end architecture behaviour;